library verilog;
use verilog.vl_types.all;
entity finaltest is
end finaltest;
