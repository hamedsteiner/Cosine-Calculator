library verilog;
use verilog.vl_types.all;
entity CosX_TB is
end CosX_TB;
